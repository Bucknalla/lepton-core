module axi_slave #(
    DATA_WIDTH = 32,
    ADDR_WIDTH = 32,
    INSTR_WIDTH = 3
)(
    input wire  S_AXI_ACLK,
    input wire  S_AXI_ARESETN,
    input wire [ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
    input wire [2 : 0] S_AXI_AWPROT,
    input wire  S_AXI_AWVALID,
    output wire  S_AXI_AWREADY,
    input wire [DATA_WIDTH-1 : 0] S_AXI_WDATA,
    input wire [(DATA_WIDTH/8)-1 : 0] S_AXI_WSTRB,
    input wire  S_AXI_WVALID,
    output wire  S_AXI_WREADY,
    output wire [1 : 0] S_AXI_BRESP,
    output wire  S_AXI_BVALID,
    input wire  S_AXI_BREADY,
    input wire [ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
    input wire [2 : 0] S_AXI_ARPROT,
    input wire  S_AXI_ARVALID,
    output wire  S_AXI_ARREADY,
    output wire [DATA_WIDTH-1 : 0] S_AXI_RDATA,
    output wire [1 : 0] S_AXI_RRESP,
    output wire  S_AXI_RVALID,
    input wire  S_AXI_RREADY,

    output wire [INSTR_WIDTH-1:0] instruction,
    output wire enable,
    
);


    
endmodule